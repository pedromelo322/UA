library ieee;
use ieee.std_logic_1164.all;

entity Controlo is
    port(
      CLOCK_50 : in std_logic;
      SW : in std_logic_vector(1 downto 0);
	  KEY : in std_logic_vector(3 downto 0);
	  LEDG : out std_logic_vector(6	downto 0);
	  LEDR : out std_logic_vector(0 downto 0);
      HEX0, HEX1, HEX2, HEX3, HEX5, HEX6, HEX7 : out std_logic_vector(6 downto 0)

    );
end Controlo;

architecture Strutural of Controlo is
    signal s_minutos0, s_minutos1, s_horas0, s_horas1 : std_logic_vector(3 downto 0) := (others => '0');
    signal s_pulse, p_pulse, minus_pulse, plus_pulse, gen_pulse, s_plus, s_minus, long_press_plus, long_press_minus: std_logic := '0';
    signal horas0, horas1, minutos0, minutos1 : std_logic_vector(6 downto 0) := (others => '0');
	signal s_set, s_modo, s_blink, blink, s_blink_h, s_blink_m, modo_ram, en_ram, OnOff: std_logic := '0';
	signal s_adress1, adress: std_logic_vector(4 downto 0) := (others => '0');
	signal s_adress0: std_logic_vector(10 downto 0) := (others => '0');
	signal s_temp, writeData: std_logic_vector(6 downto 0) := (others => '0');
	signal mux_sel : std_logic_vector(1 downto 0) := (others => '0');
	signal Tamb   : std_logic_vector(11 downto 0);
	signal tamb_dec, tamb_und, tamb_dez : std_logic_vector(3 downto 0) := (others => '0');
	signal tamb_dec_hex, tamb_und_hex, tamb_dez_hex : std_logic_vector(6 downto 0) := (others => '0');
	signal Tref : std_logic_vector(11 downto 0);

begin 


	 debounce_KEY0: entity work.DebounceUnit(Behavioral)
	
	 generic map(
		
		kHzClkFreq => 50_000,
		mSecMinInWidth => 100,
		inPolarity => '0',
		outPolarity => '1')
		
		
	 port map (
		refClk => CLOCK_50,
		dirtyIn => KEY(3),
		pulsedOut => p_pulse
	 );
		
		
	 debounce_KEY1: entity work.DebounceUnit(Behavioral)
	
	 generic map(
		
		kHzClkFreq => 50_000,
		mSecMinInWidth => 100,
		inPolarity => '0',
		outPolarity => '1')
		
		
	 port map (
		refClk => CLOCK_50,
		dirtyIn => KEY(2),
		pulsedOut => s_pulse
	 );
	 
	 debounce_KEY2: entity work.DebounceUnit(Behavioral)

	generic map(

		kHzClkFreq => 50_000,
		mSecMinInWidth => 100,
		inPolarity => '0',
		outPolarity => '1')

	
	port map (
		refClk => CLOCK_50,
		dirtyIn => KEY(1),
		pulsedOut => s_plus
	);
	
	plus_pulse <= s_plus;
	


   debounce_KEY3: entity work.DebounceUnit(Behavioral)

	generic map(

		kHzClkFreq => 50_000,
		mSecMinInWidth => 100,
		inPolarity => '0',
		outPolarity => '1')

	
	port map (
		refClk => CLOCK_50,
		dirtyIn => KEY(0),
		pulsedOut => s_minus
	);
	
	minus_pulse <= s_minus;

	 
	
	---------------------------------------------------------------------------------

	 
	controlunit_inst: entity work.ControlUnit
	  port map (
		clk              => CLOCK_50,
		set_p            => p_pulse,
		set_s            => s_pulse,
		en_7seg          => s_blink,
		modo_ram_out     => modo_ram,
		set_relogio_out  => s_set,
		modo_relogio_out => s_modo
	  );


	 
	 ---------------------------------------------------------------------------------


    pulse_generator_inst: entity work.Pulse_Generator
      port map (
        acel  => SW(1 downto 0),
        clk   => CLOCK_50,
        pulse => gen_pulse
      );

    relogio_inst: entity work.Relogio
      port map (
      en       => gen_pulse,
      clk      => CLOCK_50,
		modo 	 => s_modo,
		set 	 => s_set,
		plus 	 => plus_pulse,
		minus 	 => minus_pulse, 
		horasout => s_adress0		
      );
		
	---------------------------------------------------------------------------------
	
	RAM_inst : entity work.RAM_24_7
		port map(
			clk => CLOCK_50,
			address => adress,
			writeEnable => en_ram,
			writeData => writeData,
			readData => s_temp
		);
	
	---------------------------------------------------------------------------------

	blink_freq_inst: entity work.blink_freq
	  port map (
		clk    => CLOCK_50,
		en_in  => s_blink,
		en_out => blink
	  );

	  
	  
	blink_chs : entity work.blink_chs
		port map(
		clk => CLOCK_50,
		set => s_set,
		blink => blink,
		blink_h => s_blink_h,
		blink_m => s_blink_m
		);

	-------------------------------------------------------------------------------
		
	mux3to1_inst: entity work.mux3to1
	  port map (
		clk => CLOCK_50,
		sel => s_temp,
		y   => Tref
	  );



	controloonoff_inst: entity work.ControloOnOff
	  port map (
		clk   => CLOCK_50,
		Tref  => Tref,
		Tamb  => Tamb,
		OnOff => OnOff
	  );

	LEDR(0) <= OnOff;

	ambsimb_inst: entity work.AmbSimb
	  port map (
		clk   => gen_pulse,
		up_down => OnOff,
		counter => Tamb
	  );

	ambin_inst: entity work.AmBin
	  port map (
		clk      => CLOCK_50,
		Tamb     => Tamb,
		Tamb_dez => tamb_dez,
		Tamb_und => tamb_und,
		Tamb_dec => tamb_dec
	  );

	---------------------------------------------------------------------------------



	prog_inst: entity work.Prog
	  port map (
		en       => modo_ram,
		clk      => CLOCK_50,
		plus     => plus_pulse,
		minus    => minus_pulse,
		data_out => s_adress1
	  );

	  

	sel_inst: entity work.SEL
	  port map (
		en         => modo_ram,
		clk        => CLOCK_50,
		adress0    => s_adress0,
		adress1    => s_adress1,
		adress_out => adress,
		minutos0   => s_minutos0,
		minutos1   => s_minutos1,
		horas0     => s_horas0,
		horas1     => s_horas1
	  );


	datasel_inst: entity work.DataSEL
	  port map (
		en_ram   => en_ram,
	   data_in  => s_temp,
		modo     => modo_ram,
		clk      => CLOCK_50,
		inc      => s_pulse,
		data_out => writeData
	  );


	  
	LEDG <= writeData;

	---------------------------------------------------------------------------------
	bin7segdecoder_inst: entity work.Bin7SegDecoder
	  port map (
	   en 		=> s_blink_m,
		binInput => s_minutos0,
		decOut_n => minutos0
	  );

	bin7segdecoder_inst1: entity work.Bin7SegDecoder
	  port map (
		en 		=> s_blink_m,
		binInput => s_minutos1,
		decOut_n => minutos1
	  );	
	  
	bin7segdecoder_inst2: entity work.Bin7SegDecoder
	  port map (
	   en 		=> s_blink_h,
		binInput => s_horas0,
		decOut_n => horas0
	  );

	bin7segdecoder_inst3: entity work.Bin7SegDecoder
	  port map (
	   en 		=> s_blink_h,
		binInput => s_horas1,
		decOut_n => horas1);


	bin7segdecoder_inst4: entity work.Bin7SegDecoder
	  port map (
		en 		=> '1',
		binInput => tamb_dec,
		decOut_n => tamb_dec_hex
	  );	
	  
	bin7segdecoder_inst5: entity work.Bin7SegDecoder
	  port map (
	   en 		=> '1',
		binInput => tamb_und,
		decOut_n => tamb_und_hex
	  );

	bin7segdecoder_inst6: entity work.Bin7SegDecoder
	  port map (
	   en 		=> '1',
		binInput => tamb_dez,
		decOut_n => tamb_dez_hex);





    HEX0 <= minutos0;
    HEX1 <= minutos1;
    HEX2 <= horas0;
    HEX3 <= horas1;
	 HEX5 <= tamb_dec_hex;
    HEX6 <= tamb_und_hex;
    HEX7 <= tamb_dez_hex;

end Strutural;

